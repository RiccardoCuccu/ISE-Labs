PACKAGE constants IS
		constant N : natural := 8;
END constants;
